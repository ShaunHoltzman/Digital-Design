library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY ALUregister IS 
	PORT
		( 
			CLK                : IN STD_LOGIC;
			ALU_LD             : IN STD_LOGIC;
			ALU_OUT_EN         : IN STD_LOGIC;
			Input      			 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			ALU_OUT_FINAL      : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END ALUregister;
	
	
	ARCHITECTURE STR OF ALUregister IS 
	
	SIGNAL Data : STD_LOGIC_VECTOR(7 DOWNTO 0);
	
	BEGIN
	
		PROCESS(CLK)
	
		BEGIN
		
			IF(rising_edge(CLK)) THEN  --Synchronous load
				IF ALU_LD = '0' THEN
					Data <= Data;
				ELSIF ALU_LD = '1' THEN
					Data <= Input;
				END IF;
			END IF;
			
		END PROCESS;
		
		
		ALU_OUT_FINAL <= Data WHEN ALU_OUT_EN = '1' ELSE "ZZZZZZZZ"; --Asynchronous output enable
			
	END STR;